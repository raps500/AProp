// megafunction wizard: %Altera Multiply Adder v13.0%
// GENERATION: XML
// acog_muls.v

// Generated using ACDS version 13.0sp1 232 at 2014.04.02.21:16:19

`timescale 1 ps / 1 ps
module acog_muls (
		output wire [31:0] result,  //  result.result
		input  wire [15:0] dataa_0, // dataa_0.dataa_0
		input  wire [15:0] datab_0, // datab_0.datab_0
		input  wire        signa,   //   signa.signa
		input  wire        signb    //   signb.signb
	);

	altera_mult_add #(
		.number_of_multipliers        (1),
		.width_a                      (16),
		.width_b                      (16),
		.width_result                 (32),
		.representation_a             ("UNSIGNED"),
		.port_signa                   ("PORT_USED"),
		.signed_register_a            ("UNREGISTERED"),
		.signed_aclr_a                ("NONE"),
		.port_signb                   ("PORT_USED"),
		.representation_b             ("UNSIGNED"),
		.signed_register_b            ("UNREGISTERED"),
		.signed_aclr_b                ("NONE"),
		.output_register              ("UNREGISTERED"),
		.output_aclr                  ("NONE"),
		.multiplier1_direction        ("ADD"),
		.port_addnsub1                ("PORT_UNUSED"),
		.addnsub_multiplier_register1 ("UNREGISTERED"),
		.addnsub_multiplier_aclr1     ("NONE"),
		.multiplier3_direction        ("ADD"),
		.port_addnsub3                ("PORT_UNUSED"),
		.addnsub_multiplier_register3 ("UNREGISTERED"),
		.addnsub_multiplier_aclr3     ("NONE"),
		.input_register_a0            ("UNREGISTERED"),
		.input_register_a1            ("UNREGISTERED"),
		.input_register_a2            ("UNREGISTERED"),
		.input_register_a3            ("UNREGISTERED"),
		.input_aclr_a0                ("NONE"),
		.input_aclr_a1                ("NONE"),
		.input_aclr_a2                ("NONE"),
		.input_aclr_a3                ("NONE"),
		.input_register_b0            ("UNREGISTERED"),
		.input_register_b1            ("UNREGISTERED"),
		.input_register_b2            ("UNREGISTERED"),
		.input_register_b3            ("UNREGISTERED"),
		.input_aclr_b0                ("NONE"),
		.input_aclr_b1                ("NONE"),
		.input_aclr_b2                ("NONE"),
		.input_aclr_b3                ("NONE"),
		.scanouta_register            ("UNREGISTERED"),
		.scanouta_aclr                ("NONE"),
		.input_source_a0              ("DATAA"),
		.input_source_a1              ("DATAA"),
		.input_source_a2              ("DATAA"),
		.input_source_a3              ("DATAA"),
		.input_source_b0              ("DATAB"),
		.input_source_b1              ("DATAB"),
		.input_source_b2              ("DATAB"),
		.input_source_b3              ("DATAB"),
		.multiplier_register0         ("UNREGISTERED"),
		.multiplier_register1         ("UNREGISTERED"),
		.multiplier_register2         ("UNREGISTERED"),
		.multiplier_register3         ("UNREGISTERED"),
		.multiplier_aclr0             ("NONE"),
		.multiplier_aclr1             ("NONE"),
		.multiplier_aclr2             ("NONE"),
		.multiplier_aclr3             ("NONE"),
		.preadder_mode                ("SIMPLE"),
		.preadder_direction_0         ("ADD"),
		.preadder_direction_1         ("ADD"),
		.preadder_direction_2         ("ADD"),
		.preadder_direction_3         ("ADD"),
		.width_c                      (16),
		.input_register_c0            ("UNREGISTERED"),
		.input_register_c1            ("UNREGISTERED"),
		.input_register_c2            ("UNREGISTERED"),
		.input_register_c3            ("UNREGISTERED"),
		.input_aclr_c0                ("NONE"),
		.input_aclr_c1                ("NONE"),
		.input_aclr_c2                ("NONE"),
		.input_aclr_c3                ("NONE"),
		.width_coef                   (18),
		.coefsel0_register            ("UNREGISTERED"),
		.coefsel1_register            ("UNREGISTERED"),
		.coefsel2_register            ("UNREGISTERED"),
		.coefsel3_register            ("UNREGISTERED"),
		.coefsel0_aclr                ("NONE"),
		.coefsel1_aclr                ("NONE"),
		.coefsel2_aclr                ("NONE"),
		.coefsel3_aclr                ("NONE"),
		.coef0_0                      (0),
		.coef0_1                      (0),
		.coef0_2                      (0),
		.coef0_3                      (0),
		.coef0_4                      (0),
		.coef0_5                      (0),
		.coef0_6                      (0),
		.coef0_7                      (0),
		.coef1_0                      (0),
		.coef1_1                      (0),
		.coef1_2                      (0),
		.coef1_3                      (0),
		.coef1_4                      (0),
		.coef1_5                      (0),
		.coef1_6                      (0),
		.coef1_7                      (0),
		.coef2_0                      (0),
		.coef2_1                      (0),
		.coef2_2                      (0),
		.coef2_3                      (0),
		.coef2_4                      (0),
		.coef2_5                      (0),
		.coef2_6                      (0),
		.coef2_7                      (0),
		.coef3_0                      (0),
		.coef3_1                      (0),
		.coef3_2                      (0),
		.coef3_3                      (0),
		.coef3_4                      (0),
		.coef3_5                      (0),
		.coef3_6                      (0),
		.coef3_7                      (0),
		.accumulator                  ("NO"),
		.accum_direction              ("ADD"),
		.use_sload_accum_port         ("NO"),
		.loadconst_value              (64),
		.accum_sload_register         ("UNREGISTERED"),
		.accum_sload_aclr             ("NONE"),
		.double_accum                 ("NO"),
		.width_chainin                (1),
		.chainout_adder               ("NO"),
		.systolic_delay1              ("UNREGISTERED"),
		.systolic_aclr1               ("NONE"),
		.systolic_delay3              ("UNREGISTERED"),
		.systolic_aclr3               ("NONE"),
		.selected_device_family       ("Cyclone V")
	) acog_muls_inst (
		.result                (result),               //  result.result
		.dataa                 ({dataa_0[15:0]}),      // dataa_0.dataa_0
		.datab                 ({datab_0[15:0]}),      // datab_0.datab_0
		.signa                 (signa),                //   signa.signa
		.signb                 (signb),                //   signb.signb
		.scaninb               (16'b0000000000000000), // (terminated)
		.sourcea               (1'b0),                 // (terminated)
		.sourceb               (1'b0),                 // (terminated)
		.scanoutb              (),                     // (terminated)
		.mult01_round          (1'b0),                 // (terminated)
		.mult23_round          (1'b0),                 // (terminated)
		.mult01_saturation     (1'b0),                 // (terminated)
		.mult23_saturation     (1'b0),                 // (terminated)
		.addnsub1_round        (1'b0),                 // (terminated)
		.addnsub3_round        (1'b0),                 // (terminated)
		.mult0_is_saturated    (),                     // (terminated)
		.mult1_is_saturated    (),                     // (terminated)
		.mult2_is_saturated    (),                     // (terminated)
		.mult3_is_saturated    (),                     // (terminated)
		.output_round          (1'b0),                 // (terminated)
		.chainout_round        (1'b0),                 // (terminated)
		.output_saturate       (1'b0),                 // (terminated)
		.chainout_saturate     (1'b0),                 // (terminated)
		.chainout_sat_overflow (),                     // (terminated)
		.zero_chainout         (1'b0),                 // (terminated)
		.rotate                (1'b0),                 // (terminated)
		.shift_right           (1'b0),                 // (terminated)
		.zero_loopback         (1'b0),                 // (terminated)
		.addnsub1              (1'b1),                 // (terminated)
		.addnsub3              (1'b1),                 // (terminated)
		.clock0                (1'b1),                 // (terminated)
		.clock1                (1'b1),                 // (terminated)
		.clock2                (1'b1),                 // (terminated)
		.clock3                (1'b1),                 // (terminated)
		.ena0                  (1'b1),                 // (terminated)
		.ena1                  (1'b1),                 // (terminated)
		.ena2                  (1'b1),                 // (terminated)
		.ena3                  (1'b1),                 // (terminated)
		.aclr0                 (1'b0),                 // (terminated)
		.aclr1                 (1'b0),                 // (terminated)
		.aclr2                 (1'b0),                 // (terminated)
		.aclr3                 (1'b0),                 // (terminated)
		.scanina               (16'b0000000000000000), // (terminated)
		.scanouta              (),                     // (terminated)
		.coefsel0              (3'b000),               // (terminated)
		.coefsel1              (3'b000),               // (terminated)
		.coefsel2              (3'b000),               // (terminated)
		.coefsel3              (3'b000),               // (terminated)
		.datac                 (16'b0000000000000000), // (terminated)
		.accum_sload           (1'b0),                 // (terminated)
		.sload_accum           (1'b0),                 // (terminated)
		.chainin               (1'b0)                  // (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2014 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_mult_add" version="13.0" >
// Retrieval info: 	<generic name="number_of_multipliers" value="1" />
// Retrieval info: 	<generic name="width_a" value="16" />
// Retrieval info: 	<generic name="width_b" value="16" />
// Retrieval info: 	<generic name="width_result" value="32" />
// Retrieval info: 	<generic name="gui_4th_asynchronous_clear" value="false" />
// Retrieval info: 	<generic name="gui_associated_clock_enable" value="false" />
// Retrieval info: 	<generic name="gui_representation_a" value="VARIABLE" />
// Retrieval info: 	<generic name="gui_register_signa" value="false" />
// Retrieval info: 	<generic name="gui_register_signa_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_register_signa_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_representation_b" value="VARIABLE" />
// Retrieval info: 	<generic name="gui_register_signb" value="false" />
// Retrieval info: 	<generic name="gui_register_signb_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_register_signb_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_a_shiftout" value="false" />
// Retrieval info: 	<generic name="gui_b_shiftout" value="false" />
// Retrieval info: 	<generic name="gui_output_register" value="false" />
// Retrieval info: 	<generic name="gui_output_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_output_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_multiplier1_direction" value="ADD" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_register1" value="false" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_register1_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_aclr1" value="NONE" />
// Retrieval info: 	<generic name="gui_multiplier3_direction" value="ADD" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_register3" value="false" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_register3_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_addnsub_multiplier_aclr3" value="NONE" />
// Retrieval info: 	<generic name="gui_input_register_a" value="false" />
// Retrieval info: 	<generic name="gui_input_register_a_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_input_register_a_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_input_register_b" value="false" />
// Retrieval info: 	<generic name="gui_input_register_b_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_input_register_b_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_multiplier_a_input" value="Multiplier input" />
// Retrieval info: 	<generic name="gui_scanouta_register" value="false" />
// Retrieval info: 	<generic name="gui_scanouta_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_scanouta_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_multiplier_b_input" value="Multiplier input" />
// Retrieval info: 	<generic name="gui_multiplier_register" value="false" />
// Retrieval info: 	<generic name="gui_multiplier_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_multiplier_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="preadder_mode" value="SIMPLE" />
// Retrieval info: 	<generic name="gui_preadder_direction" value="ADD" />
// Retrieval info: 	<generic name="width_c" value="16" />
// Retrieval info: 	<generic name="gui_datac_input_register" value="false" />
// Retrieval info: 	<generic name="gui_datac_input_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_datac_input_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="width_coef" value="18" />
// Retrieval info: 	<generic name="gui_coef_register" value="false" />
// Retrieval info: 	<generic name="gui_coef_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_coef_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="coef0_0" value="0" />
// Retrieval info: 	<generic name="coef0_1" value="0" />
// Retrieval info: 	<generic name="coef0_2" value="0" />
// Retrieval info: 	<generic name="coef0_3" value="0" />
// Retrieval info: 	<generic name="coef0_4" value="0" />
// Retrieval info: 	<generic name="coef0_5" value="0" />
// Retrieval info: 	<generic name="coef0_6" value="0" />
// Retrieval info: 	<generic name="coef0_7" value="0" />
// Retrieval info: 	<generic name="coef1_0" value="0" />
// Retrieval info: 	<generic name="coef1_1" value="0" />
// Retrieval info: 	<generic name="coef1_2" value="0" />
// Retrieval info: 	<generic name="coef1_3" value="0" />
// Retrieval info: 	<generic name="coef1_4" value="0" />
// Retrieval info: 	<generic name="coef1_5" value="0" />
// Retrieval info: 	<generic name="coef1_6" value="0" />
// Retrieval info: 	<generic name="coef1_7" value="0" />
// Retrieval info: 	<generic name="coef2_0" value="0" />
// Retrieval info: 	<generic name="coef2_1" value="0" />
// Retrieval info: 	<generic name="coef2_2" value="0" />
// Retrieval info: 	<generic name="coef2_3" value="0" />
// Retrieval info: 	<generic name="coef2_4" value="0" />
// Retrieval info: 	<generic name="coef2_5" value="0" />
// Retrieval info: 	<generic name="coef2_6" value="0" />
// Retrieval info: 	<generic name="coef2_7" value="0" />
// Retrieval info: 	<generic name="coef3_0" value="0" />
// Retrieval info: 	<generic name="coef3_1" value="0" />
// Retrieval info: 	<generic name="coef3_2" value="0" />
// Retrieval info: 	<generic name="coef3_3" value="0" />
// Retrieval info: 	<generic name="coef3_4" value="0" />
// Retrieval info: 	<generic name="coef3_5" value="0" />
// Retrieval info: 	<generic name="coef3_6" value="0" />
// Retrieval info: 	<generic name="coef3_7" value="0" />
// Retrieval info: 	<generic name="accumulator" value="NO" />
// Retrieval info: 	<generic name="accum_direction" value="ADD" />
// Retrieval info: 	<generic name="gui_ena_preload_const" value="false" />
// Retrieval info: 	<generic name="gui_accumulate_port_select" value="0" />
// Retrieval info: 	<generic name="loadconst_value" value="64" />
// Retrieval info: 	<generic name="gui_accum_sload_register_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_accum_sload_register_aclr" value="NONE" />
// Retrieval info: 	<generic name="gui_double_accum" value="false" />
// Retrieval info: 	<generic name="gui_chainout_adder" value="false" />
// Retrieval info: 	<generic name="chainout_adder" value="NO" />
// Retrieval info: 	<generic name="gui_systolic_delay" value="false" />
// Retrieval info: 	<generic name="gui_systolic_delay_clock" value="CLOCK0" />
// Retrieval info: 	<generic name="gui_systolic_delay_aclr" value="NONE" />
// Retrieval info: 	<generic name="selected_device_family" value="Cyclone V" />
// Retrieval info: 	<generic name="reg_autovec_sim" value="false" />
// Retrieval info: </instance>
// IPFS_FILES : acog_muls.vo
// RELATED_FILES: acog_muls.v
