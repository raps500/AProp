/*
 * Testbench for the alu
 *
 */

`include "acog_alu.v"
module tb_alu();

reg clk, C, Z;
reg [31:0] S, D;
reg [8:0] pc_plus_1;
reg [5:0] opcode;
wire [31:0] alu_q;
wire alu_c;
wire alu_z;


acog_alu alu(
	.clk_in(clk),
	.opcode_in(opcode),
	.flag_c_in(C),
	.flag_z_in(Z),
	.s_in(S),
	.s_negative_in(32'h0-S),
	.d_in(D),
	.pc_plus_1_in(pc_plus_1),
	.d_is_zero_in(D == 32'h0),
	.flag_c_o(alu_c),
	.flag_z_o(alu_z),
	.q_o(alu_q)
	);
	
initial
	begin
	$dumpfile("tb_alu.vcd");
	$dumpvars(0, tb_alu);
	$display("ROR     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ROR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ROL     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ROL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SHR     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SHR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SHL     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SHL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("RCR     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_RCR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("RCL     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_RCL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SAR     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SAR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("REV     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_REV;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MINS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MINS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MAXS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MAXS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MIN     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MIN	;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MAX     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MAX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MOVS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MOVS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MOVD    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MOVD;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MOVI    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MOVI;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("JMPRET  ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_JMPRET;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("AND     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_AND;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ANDN    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ANDN;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("OR      ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_OR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("XOR     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_XOR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MUXC    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MUXC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MUXNC   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MUXNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MUXNZ   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MUXNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MUXZ    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MUXZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ADD     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ADD;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUB     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUB;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ADDABS  ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ADDABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUBABS  ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUBABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUMC    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUMC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUMNC   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUMNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUMZ    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUMZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUMNZ   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUMNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("MOV     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_MOV;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("NEG     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_NEG;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ABS     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ABSNEG  ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ABSNEG;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("NEGC    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_NEGC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("NEGZ    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_NEGZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("NEGNC   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_NEGNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("NEGNZ   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_NEGNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("CMPS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_CMPS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("CMPSX   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_CMPSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ADDX    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ADDX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUBX    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUBX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ADDS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ADDS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUBS    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUBS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("ADDSX   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_ADDSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("SUBSX   ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_SUBSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("CMPSUB  ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_CMPSUB;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("DJNZ    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_DJNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("TJNZ    ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_TJNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("TJZ     ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_TJZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("WAITPEQ ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_WAITPEQ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("WAITPNE ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_WAITPNE;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("WAITCNT ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_WAITCNT;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	$display("WAITVID ---D---- ---S---- ZC = ---Q---- ZC");

	#1
    opcode = `I_WAITVID;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("        %08x %08x %1x%1x = %08x %1x%1x", D, S, Z, C, alu_q, alu_z, alu_c);
    end
endmodule
