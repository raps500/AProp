/*
 * Testbench for the alu
 *
 */

`include "acog_alu.v"
module tb_alu();

reg clk, C, Z;
reg [31:0] S, D;
reg [8:0] pc_plus_1;
reg [5:0] opcode;
wire [31:0] alu_q;
wire alu_c;
wire alu_z;


acog_alu alu(
	.clk_in(clk),
	.opcode_in({opcode, 26'h0 }),
	.flag_c_in(C),
	.flag_z_in(Z),
	.s_in(S),
	.d_in(D),
	.pc_plus_1_in(pc_plus_1),
	.flag_c_o(alu_c),
	.flag_z_o(alu_z),
	.q_o(alu_q)
	);
	
initial
	begin
	$dumpfile("tb_alu.vcd");
	$dumpvars(0, tb_alu);
	$display("ROR   ---Q---- CZ");

	#1
    opcode = `I_ROR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ROL   ---Q---- CZ");

	#1
    opcode = `I_ROL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SHR   ---Q---- CZ");

	#1
    opcode = `I_SHR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SHL   ---Q---- CZ");

	#1
    opcode = `I_SHL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("RCR   ---Q---- CZ");

	#1
    opcode = `I_RCR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("RCL   ---Q---- CZ");

	#1
    opcode = `I_RCL;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SAR   ---Q---- CZ");

	#1
    opcode = `I_SAR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("REV   ---Q---- CZ");

	#1
    opcode = `I_REV;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MINS  ---Q---- CZ");

	#1
    opcode = `I_MINS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MAXS  ---Q---- CZ");

	#1
    opcode = `I_MAXS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MIN   ---Q---- CZ");

	#1
    opcode = `I_MIN	;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MAX   ---Q---- CZ");

	#1
    opcode = `I_MAX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MOVS  ---Q---- CZ");

	#1
    opcode = `I_MOVS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MOVD  ---Q---- CZ");

	#1
    opcode = `I_MOVD;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MOVI  ---Q---- CZ");

	#1
    opcode = `I_MOVI;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("JMPRET---Q---- CZ");

	#1
    opcode = `I_JMPRET;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("AND   ---Q---- CZ");

	#1
    opcode = `I_AND;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ANDN  ---Q---- CZ");

	#1
    opcode = `I_ANDN;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("OR    ---Q---- CZ");

	#1
    opcode = `I_OR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("XOR   ---Q---- CZ");

	#1
    opcode = `I_XOR;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MUXC  ---Q---- CZ");

	#1
    opcode = `I_MUXC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MUXNC ---Q---- CZ");

	#1
    opcode = `I_MUXNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MUXNZ ---Q---- CZ");

	#1
    opcode = `I_MUXNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MUXZ  ---Q---- CZ");

	#1
    opcode = `I_MUXZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ADD   ---Q---- CZ");

	#1
    opcode = `I_ADD;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUB   ---Q---- CZ");

	#1
    opcode = `I_SUB;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ADDABS---Q---- CZ");

	#1
    opcode = `I_ADDABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUBABS---Q---- CZ");

	#1
    opcode = `I_SUBABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUMC  ---Q---- CZ");

	#1
    opcode = `I_SUMC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUMNC ---Q---- CZ");

	#1
    opcode = `I_SUMNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUMZ  ---Q---- CZ");

	#1
    opcode = `I_SUMZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUMNZ ---Q---- CZ");

	#1
    opcode = `I_SUMNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("MOV   ---Q---- CZ");

	#1
    opcode = `I_MOV;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("NEG   ---Q---- CZ");

	#1
    opcode = `I_NEG;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ABS   ---Q---- CZ");

	#1
    opcode = `I_ABS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ABSNEG---Q---- CZ");

	#1
    opcode = `I_ABSNEG;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("NEGC  ---Q---- CZ");

	#1
    opcode = `I_NEGC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("NEGZ  ---Q---- CZ");

	#1
    opcode = `I_NEGZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("NEGNC ---Q---- CZ");

	#1
    opcode = `I_NEGNC;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("NEGNZ ---Q---- CZ");

	#1
    opcode = `I_NEGNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("CMPS  ---Q---- CZ");

	#1
    opcode = `I_CMPS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("CMPSX ---Q---- CZ");

	#1
    opcode = `I_CMPSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ADDX  ---Q---- CZ");

	#1
    opcode = `I_ADDX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUBX  ---Q---- CZ");

	#1
    opcode = `I_SUBX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ADDS  ---Q---- CZ");

	#1
    opcode = `I_ADDS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUBS  ---Q---- CZ");

	#1
    opcode = `I_SUBS;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("ADDSX ---Q---- CZ");

	#1
    opcode = `I_ADDSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("SUBSX ---Q---- CZ");

	#1
    opcode = `I_SUBSX;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("CMPSUB---Q---- CZ");

	#1
    opcode = `I_CMPSUB;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("DJNZ  ---Q---- CZ");

	#1
    opcode = `I_DJNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("TJNZ  ---Q---- CZ");

	#1
    opcode = `I_TJNZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("TJZ   ---Q---- CZ");

	#1
    opcode = `I_TJZ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("WAITPEQ---Q---- CZ");

	#1
    opcode = `I_WAITPEQ;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("WAITPNE---Q---- CZ");

	#1
    opcode = `I_WAITPNE;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("WAITCNT---Q---- CZ");

	#1
    opcode = `I_WAITCNT;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	$display("WAITVID---Q---- CZ");

	#1
    opcode = `I_WAITVID;
	S = 32'h00000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("00 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("01 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("02 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("03 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("04 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("05 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("06 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("07 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("08 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("09 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("0c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("0d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("0e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("0f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("10 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("11 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("12 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("13 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("14 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("15 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("16 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("17 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("18 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("19 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("1c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("1d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("1e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("1f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("20 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("21 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("22 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("23 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("24 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("25 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("26 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("27 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("28 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("29 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("2c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("2d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("2e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("2f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("30 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("31 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("32 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("33 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("34 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("35 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("36 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("37 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("38 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("39 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("3c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("3d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("3e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("3f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("40 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("41 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("42 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("43 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("44 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("45 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("46 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("47 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("48 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("49 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("4c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("4d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("4e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("4f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("50 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("51 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("52 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("53 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("54 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("55 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("56 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("57 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("58 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("59 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h00000002;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("5c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("5d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("5e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("5f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("60 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("61 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("62 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("63 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("64 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("65 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("66 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("67 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("68 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("69 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("6c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("6d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("6e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("6f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("70 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("71 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("72 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("73 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("74 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("75 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("76 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("77 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("78 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("79 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h7fffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("7c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("7d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("7e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("7f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("80 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("81 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("82 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("83 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("84 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("85 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("86 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("87 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("88 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("89 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("8c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("8d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("8e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("8f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("90 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("91 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("92 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("93 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("94 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("95 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("96 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("97 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("98 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("99 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9a %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9b %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000000;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("9c %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("9d %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("9e %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("9f %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("a6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("a7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("a8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("a9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("aa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ab %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ac %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ad %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ae %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("af %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("b6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("b7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("b8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("b9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ba %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'h80000001;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("bc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("bd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("be %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("bf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("c6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("c7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("c8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("c9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ca %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("cc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("cd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ce %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("cf %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("d6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("d7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("d8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("d9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("da %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("db %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hfffffffe;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("dc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("dd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("de %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("df %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("e6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("e7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h00000002;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("e8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("e9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ea %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("eb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h7fffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("ec %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("ed %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("ee %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ef %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000000;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f0 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f1 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f2 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f3 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'h80000001;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f4 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f5 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("f6 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("f7 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hfffffffe;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("f8 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("f9 %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fa %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("fb %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	S = 32'hffffffff;
	D = 32'hffffffff;
	C = 1'b0;
	Z = 1'b0;
	#1 $display("fc %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b0;
	#1 $display("fd %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b0;
	Z = 1'b1;
	#1 $display("fe %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
	#1
	C = 1'b1;
	Z = 1'b1;
	#1 $display("ff %02x %08x %1x%1x", opcode, alu_q, alu_c, alu_z);
    end
endmodule
