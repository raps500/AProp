/* 
 * ACog - Fetch unit
 *
 * 
 */
`include "acog_defs.v" 

module acog_if(
	input wire clk_in,
	input wire [1:0] state_in
	);
	


	
endmodule
